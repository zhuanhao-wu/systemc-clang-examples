module sreg_0(
input wire [0:0] clk,
input wire [0:0] reset 
);


always @(*) begin: mc_io

reg m_port;
reg s_port;
reg s_port;
end // mc_io
endmodule // sreg_0
module sreg_1(
input wire [0:0] clk,
input wire [0:0] reset 
);


always @(*) begin: mc_io

reg m_port;
reg s_port;
reg s_port;
end // mc_io
endmodule // sreg_1
module sreg_2(
input wire [0:0] clk,
input wire [0:0] reset 
);


always @(*) begin: mc_io

reg m_port;
reg s_port;
reg s_port;
end // mc_io
endmodule // sreg_2
module test_0(
 
);


always @(*) begin: mc_test


end // mc_test
endmodule // test_0