module fa_0(
input wire [0:0] a,
input wire [0:0] b,
input wire [0:0] cin,
output reg [0:0] cout,
output reg [0:0] s 
);



endmodule // fa_0
module fa_1(
input wire [0:0] a,
input wire [0:0] b,
input wire [0:0] cin,
output reg [0:0] cout,
output reg [0:0] s 
);



endmodule // fa_1
module fa_2(
input wire [0:0] a,
input wire [0:0] b,
input wire [0:0] cin,
output reg [0:0] cout,
output reg [0:0] s 
);



endmodule // fa_2
module fa_3(
input wire [0:0] a,
input wire [0:0] b,
input wire [0:0] cin,
output reg [0:0] cout,
output reg [0:0] s 
);



endmodule // fa_3