module top_0(
input wire clk,
input wire integer in_port,
output reg integer out_port 
);
sc_event aev;
integer v;
integer w;
integer x;
integer y;


endmodule // top_0
module top_1(
input wire clk,
input wire integer in_port,
output reg integer out_port 
);
sc_event aev;
integer v;
integer w;
integer x;
integer y;


endmodule // top_1