module top_0(
input wire clk,
input wire integer int_port 
);
integer var;
integer x;
integer y;


endmodule // top_0