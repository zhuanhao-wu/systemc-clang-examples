module top_0(
input wire clk,
input wire integer in_port,
output reg integer out_port 
);
integer var;
integer x;
integer y;


endmodule // top_0