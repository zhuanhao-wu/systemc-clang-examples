module producer_0(
input wire [0:0] clock,
input wire integer in1,
output reg integer out,
output reg [0:0] ready 
);



endmodule // producer_0